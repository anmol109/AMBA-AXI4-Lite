module AXI_lite();